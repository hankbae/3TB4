module Ass2(
	input CLOCK,
			n_R_W,
			request,
			ack,
	input [3:0] address_master,
					addressBuff_slave,
					data_master,
	input [3:0] data_slave,
	input [7:0] dataBuff_master,
	output rand
	);
endmodule 