
module lab2tut (input CLOCK_50,
					input [2:0] KEY,
					output [6:0] HEX0,
					HEX1,
					HEX2,
					HEX3,
					HEX4,
					HEX5);
					
always @(posedge CLOCK_50)
begin
		


end
					
					
					
					
endmodule
